module ALU (output[7:0] reg_out, output[7:0] SREG, input[2:0] function_select_lines, input[7:0] operandA, input[7:0] operandB);

endmodule // ALU
