module dataMemory (input clk);

endmodule
