module CU (input[32:0] instruction);
    wire[7:0] operandA, operandB;
    wire[4:0] opcode;

    
endmodule
