module cache (input[])
