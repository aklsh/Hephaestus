module EU ();
    
endmodule
